
module toplevel(CLOCK_50, SW, KEY, AUD_ADCDAT,

	// Bidirectionals
	AUD_BCLK,
	AUD_ADCLRCK,
	AUD_DACLRCK,

	FPGA_I2C_SDAT,

	// Outputs
	AUD_XCK,
	AUD_DACDAT,

	FPGA_I2C_SCLK, song_data);

	input CLOCK_50;
	input [3:0] SW;
	input [0:0] KEY;

	wire [7:0] memory_address_song;
	wire [31:0] song_data_out;
	output [31:0] song_data;

	
	//song_data = song_data_out;
	
	//inputs
	input				AUD_ADCDAT;

	// Bidirectionals
	inout				AUD_BCLK;
	inout				AUD_ADCLRCK;
	inout				AUD_DACLRCK;

	inout				FPGA_I2C_SDAT;

	// Outputs
	output				AUD_XCK;
	output				AUD_DACDAT;

	output				FPGA_I2C_SCLK;
	
	//internal wires: 
	wire				audio_in_available;
	wire		[31:0]	left_channel_audio_in;
	wire		[31:0]	right_channel_audio_in;
	wire				read_audio_in;

	wire				audio_out_allowed;
	wire		[31:0]	left_channel_audio_out;
	wire		[31:0]	right_channel_audio_out;
	wire				write_audio_out;
	
	//Internal Registers: 
	//reg [10:0] delay_cnt;
	//wire [10:0] delay;

	//reg snd;
	
	//counter
//	always @(posedge CLOCK_50)
//	if(delay_cnt == delay) begin
//		delay_cnt <= 0;
//		snd <= !snd; //pulse
//	end else delay_cnt <= delay_cnt + 1;
//assign delay = 11'd1042; //constant audio output/ 
/*****************************************************************************
 *                            Combinational Logic                            *
 *****************************************************************************/
 
	reg [15:0] address;
	reg [15:0] counter;
	//audio_out_allowed is technically the enable signal
	
	//values to set to one: 
	//assign write_audio_out = 1'b1;
	
	always @(posedge CLOCK_50) begin
		if(~KEY[0]) begin
		address <= 16'd0;
		counter <= 16'd0;
		end
		if (audio_out_allowed) begin
			address <= counter; 
			counter <= counter + 16'd1;
		end
	  if (counter == 16'd45852) counter <= 16'd0;	
	  if (audio_out_allowed == 0) begin
	  counter <= counter + 16'd0; //extra safety
	  address <= address + 16'd0; //does nothing.
	  end
	end
	
	//reads address bit by bit
	ram32x4 r1(.address(address), .clock(CLOCK_50), .data(32'b0), .wren(1'b0), .q(song_data_out)); //enables read - only.
	
	assign left_channel_audio_out	= song_data_out;
	assign right_channel_audio_out = song_data_out;
		
	assign read_audio_in			= audio_in_available & audio_out_allowed;
	assign write_audio_out			= audio_in_available & audio_out_allowed;

	
	//fuck my ass setting these to 0.
//	assign read_audio_in = 1'b0;
//	assign audio_in_available = 1'b0;
//	assign left_channel_audio_in = 1'b0;
//	assign right_channel_audio_in = 1'b0;

	
	Audio_Controller Audio_Controller (
	// Inputs
	.CLOCK_50						(CLOCK_50),
	.reset						(~KEY[0]),

	.clear_audio_in_memory		(),
	.read_audio_in				(read_audio_in),
	
	.clear_audio_out_memory		(),
	.left_channel_audio_out		(left_channel_audio_out),
	.right_channel_audio_out	(right_channel_audio_out),
	.write_audio_out			(write_audio_out),

	.AUD_ADCDAT					(AUD_ADCDAT),

	// Bidirectionals
	.AUD_BCLK					(AUD_BCLK),
	.AUD_ADCLRCK				(AUD_ADCLRCK),
	.AUD_DACLRCK				(AUD_DACLRCK),


	// Outputs
	.audio_in_available			(audio_in_available),
	.left_channel_audio_in		(left_channel_audio_in),
	.right_channel_audio_in		(right_channel_audio_in),

	.audio_out_allowed			(audio_out_allowed),

	.AUD_XCK					(AUD_XCK),
	.AUD_DACDAT					(AUD_DACDAT)

);

endmodule

//old code 
//assign read_audio_in	= snd? audio_in_available & audio_out_allowed : 0;
//assign write_audio_out			= audio_in_available & audio_out_allowed;

	//assign write_audio_out = 0;
	//assign audio_out_allowed = 1'b1;
	
	//assign audio_read_in = 1'b1;
	
	//assign left_channel_audio_in; //nani
	//assign right_channel_audio_in;
	//assign read_audio_in = 1'b1; //pulse this

	
//module ram32x4 (
//	address,
//	clock,
//	data,
//	wren,
//	q);
//endmodule

//module audiotest (
//	// Inputs
//	CLOCK_50,
//	KEY,
//
//	AUD_ADCDAT,
//
//	// Bidirectionals
//	AUD_BCLK,
//	AUD_ADCLRCK,
//	AUD_DACLRCK,
//
//	FPGA_I2C_SDAT,
//
//	// Outputs
//	AUD_XCK,
//	AUD_DACDAT,
//
//	FPGA_I2C_SCLK,
//	//SW
//);
//
///*****************************************************************************
// *                           Parameter Declarations                          *
// *****************************************************************************/
//
//
///*****************************************************************************
// *                             Port Declarations                             *
// *****************************************************************************/
//// Inputs
//input				CLOCK_50;
//input		[3:0]	KEY;
//input		[3:0]	SW;
//
//input				AUD_ADCDAT;
//
//// Bidirectionals
//inout				AUD_BCLK;
//inout				AUD_ADCLRCK;
//inout				AUD_DACLRCK;
//
//inout				FPGA_I2C_SDAT;
//
//// Outputs
//output				AUD_XCK;
//output				AUD_DACDAT;
//
//output				FPGA_I2C_SCLK;
//
///*****************************************************************************
// *                 Internal Wires and Registers Declarations                 *
// *****************************************************************************/
//// Internal Wires
//wire				audio_in_available;
//wire		[31:0]	left_channel_audio_in;
//wire		[31:0]	right_channel_audio_in;
//wire				read_audio_in;
//
//wire				audio_out_allowed;
//wire		[31:0]	left_channel_audio_out;
//wire		[31:0]	right_channel_audio_out;
//wire				write_audio_out;
//
//// Internal Registers
//
//reg [18:0] delay_cnt;
//wire [18:0] delay;
//
//reg snd;
//
//// State Machine Registers
//
///*****************************************************************************
// *                         Finite State Machine(s)                           *
// *****************************************************************************/
//
//
///*****************************************************************************
// *                             Sequential Logic                              *
// *****************************************************************************/
//
//always @(posedge CLOCK_50)
//	if(delay_cnt == delay) begin
//		delay_cnt <= 0;
//		snd <= !snd;
//	end else delay_cnt <= delay_cnt + 1;
//
///*****************************************************************************
// *                            Combinational Logic                            *
// *****************************************************************************/
//
//assign delay = {SW[3:0], 15'd3000};
//
//wire [31:0] sound = (SW == 0) ? 0 : snd ? 32'd10000000 : -32'd10000000;
//
//
//assign read_audio_in			= audio_in_available & audio_out_allowed;
//
//assign left_channel_audio_out	= left_channel_audio_in+sound;
//assign right_channel_audio_out	= right_channel_audio_in+sound;
//assign write_audio_out			= audio_in_available & audio_out_allowed;
//
///*****************************************************************************
// *                              Internal Modules                             *
// *****************************************************************************/
//
//Audio_Controller Audio_Controller (
//	// Inputs
//	.CLOCK_50						(CLOCK_50),
//	.reset						(~KEY[0]),
//
//	.clear_audio_in_memory		(),
//	.read_audio_in				(read_audio_in),
//	
//	.clear_audio_out_memory		(),
//	.left_channel_audio_out		(left_channel_audio_out),
//	.right_channel_audio_out	(right_channel_audio_out),
//	.write_audio_out			(write_audio_out),
//
//	.AUD_ADCDAT					(AUD_ADCDAT),
//
//	// Bidirectionals
//	.AUD_BCLK					(AUD_BCLK),
//	.AUD_ADCLRCK				(AUD_ADCLRCK),
//	.AUD_DACLRCK				(AUD_DACLRCK),
//
//
//	// Outputs
//	.audio_in_available			(audio_in_available),
//	.left_channel_audio_in		(left_channel_audio_in),
//	.right_channel_audio_in		(right_channel_audio_in),
//
//	.audio_out_allowed			(audio_out_allowed),
//
//	.AUD_XCK					(AUD_XCK),
//	.AUD_DACDAT					(AUD_DACDAT)
//
//);
//
//avconf #(.USE_MIC_INPUT(1)) avc (
//	.FPGA_I2C_SCLK					(FPGA_I2C_SCLK),
//	.FPGA_I2C_SDAT					(FPGA_I2C_SDAT),
//	.CLOCK_50					(CLOCK_50),
//	.reset						(~KEY[0])
//);
//
//endmodule

