
module DE1_SoC_Audio_Example (
	// Inputs
	CLOCK_50,
	KEY, HEX0,HEX1, HEX2, HEX3, HEX4, HEX5,

	AUD_ADCDAT,

	// Bidirectionals
	AUD_BCLK,
	AUD_ADCLRCK,
	AUD_DACLRCK,

	FPGA_I2C_SDAT,

	// Outputs
	AUD_XCK,
	AUD_DACDAT,

	FPGA_I2C_SCLK,
	SW
);

/*****************************************************************************
 *                           Parameter Declarations                          *
 *****************************************************************************/


/*****************************************************************************
 *                             Port Declarations                             *
 *****************************************************************************/
// Inputs
input				CLOCK_50;
input		[3:0]	KEY;
input		[3:0]	SW;

input				AUD_ADCDAT;

// Bidirectionals
inout				AUD_BCLK;
inout				AUD_ADCLRCK;
inout				AUD_DACLRCK;

inout				FPGA_I2C_SDAT;

// Outputs
output				AUD_XCK;
output				AUD_DACDAT;

output				FPGA_I2C_SCLK;
output [6:0] HEX0 , HEX1, HEX2, HEX3, HEX4, HEX5;

/*****************************************************************************
 *                 Internal Wires and Registers Declarations                 *
 *****************************************************************************/
// Internal Wires
wire				audio_in_available;
wire		[31:0]	left_channel_audio_in;
wire		[31:0]	right_channel_audio_in;
wire				read_audio_in;

wire				audio_out_allowed;
wire		[31:0]	left_channel_audio_out;
wire		[31:0]	right_channel_audio_out;
wire				write_audio_out;

// Internal Registers

//reg [18:0] delay_cnt;
//wire [18:0] delay;
reg [18:0] delay_cnt;
wire [18:0] delay;


reg [18:0] delay_cnt2;
wire [18:0] delay2;

reg snd;

reg [15:0] freq2;
wire [19:0] audio_out; // output of the ram
reg [26:0] frequency_counter;
reg [9:0] address;
wire reset = ~KEY[0];

testram test(.address(address), .clock(CLOCK_50), .data(18'b0), .wren(1'b0), .q(audio_out)); 
hex_decoder h1(.hex_digit(address [3:0]), .segments(HEX0));
hex_decoder h2(.hex_digit(address [7:4]), .segments(HEX1));
hex_decoder h3(.hex_digit({2'b0, audio_out [9:8]}), .segments(HEX2));
//hex_decoder h4(.hex_digit(audio_out [15:12]), .segments(HEX3));
//hex_decoder h5(.hex_digit({2'b0, audio_out [17:16]}), .segments(HEX4));
//hex_decoder h6(.hex_digit(3'd4), .segments(HEX5));

// State Machine Registers

/*****************************************************************************
 *                         Finite State Machine(s)                           *
 *****************************************************************************/


/*****************************************************************************
 *                             Sequential Logic                              *
 *****************************************************************************/
//change this value 
reg [20:0] mif_lines = 10'd252;
reg [26:0] limit = 27'd9200000;
reg [20:0] tempo_change_one = 10'd197;

always @(posedge CLOCK_50)
		if(delay_cnt == delay) begin
			delay_cnt <= 0;
			snd <= !snd;
		end else delay_cnt <= delay_cnt + 1;

// rate divider
always @(posedge CLOCK_50) begin
		if (reset) address <= 0;
		if (frequency_counter == limit) begin 
			frequency_counter <= 27'b0;
			if (address == mif_lines) begin
				address <= 0;
				limit <= 27'd9200000;
			end
			if (address < mif_lines)
				address <= address + 1;
			if (address == tempo_change_one) //speeding the tempo up.
			   limit <= 27'd7800000;
			end
		else 
			frequency_counter <= frequency_counter + 1;
	end

/*****************************************************************************
 *                            Combinational Logic                            *
 *****************************************************************************/

assign delay = audio_out;

wire [31:0] sound = (SW == 0) ? 0 : snd ? 32'd1000000000 : -32'd1000000000;


assign read_audio_in			= audio_in_available & audio_out_allowed;

assign left_channel_audio_out	= left_channel_audio_in+sound;
assign right_channel_audio_out	= right_channel_audio_in+sound;
assign write_audio_out			= audio_in_available & audio_out_allowed;

/*****************************************************************************
 *                              Internal Modules                             *
 *****************************************************************************/

Audio_Controller Audio_Controller (
	// Inputs
	.CLOCK_50						(CLOCK_50),
	.reset						(~KEY[0]),

	.clear_audio_in_memory		(),
	.read_audio_in				(read_audio_in),
	
	.clear_audio_out_memory		(),
	.left_channel_audio_out		(left_channel_audio_out),
	.right_channel_audio_out	(right_channel_audio_out),
	.write_audio_out			(write_audio_out),

	.AUD_ADCDAT					(AUD_ADCDAT),

	// Bidirectionals
	.AUD_BCLK					(AUD_BCLK),
	.AUD_ADCLRCK				(AUD_ADCLRCK),
	.AUD_DACLRCK				(AUD_DACLRCK),


	// Outputs
	.audio_in_available			(audio_in_available),
	.left_channel_audio_in		(left_channel_audio_in),
	.right_channel_audio_in		(right_channel_audio_in),

	.audio_out_allowed			(audio_out_allowed),

	.AUD_XCK					(AUD_XCK),
	.AUD_DACDAT					(AUD_DACDAT)

);

avconf #(.USE_MIC_INPUT(1)) avc (
	.FPGA_I2C_SCLK					(FPGA_I2C_SCLK),
	.FPGA_I2C_SDAT					(FPGA_I2C_SDAT),
	.CLOCK_50					(CLOCK_50),
	.reset						(~KEY[0])
);

endmodule

module hex_decoder(hex_digit, segments);
    input [3:0] hex_digit;
    output reg [6:0] segments;
   
    always @(*)
        case (hex_digit)
            4'h0: segments = 7'b100_0000;
            4'h1: segments = 7'b111_1001;
            4'h2: segments = 7'b010_0100;
            4'h3: segments = 7'b011_0000;
            4'h4: segments = 7'b001_1001;
            4'h5: segments = 7'b001_0010;
            4'h6: segments = 7'b000_0010;
            4'h7: segments = 7'b111_1000;
            4'h8: segments = 7'b000_0000;
            4'h9: segments = 7'b001_1000;
            4'hA: segments = 7'b000_1000;
            4'hB: segments = 7'b000_0011;
            4'hC: segments = 7'b100_0110;
            4'hD: segments = 7'b010_0001;
            4'hE: segments = 7'b000_0110;
            4'hF: segments = 7'b000_1110;   
            default: segments = 7'h7f;
        endcase
endmodule

